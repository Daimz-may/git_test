module test(
a,b,c);
input [3:0] a;
input [3:0] b;
output [4:0] c;

c=a+b;
	
endmodule
